import params::*;
import typesPkg::*;

module mii_module (
    input logic clk, // main clock
    input logic eth_txck_in, // internal transmit clock 125 MHz -1GBit / 25MHz - 100Mbit
    input logic eth_txclk_phy, // transmit clock from a pll to the mii interface 125 MHz -1GBit / 25MHz - 100Mbit
    input logic rst_n, // hold in reset state before all the initialization is done

    input logic eth_rxclk, // clock generated by the mii rx interface 125 MHz -1GBit / 25MHz - 100Mbit
    input logic eth_rxdv,
    input logic [3:0] eth_rxd,
    output logic eth_txclk,
    output logic eth_txdv,
    output logic [3:0] eth_txd,

    output logic valid_rx,      /* Valid data, strobe after preamble including crc */
    output logic [7:0] data_rx, /* RX data */

    input mii_tx_t mii_tx, // tx stream from queue

    output mii_rx_status_t rx_stat,
    input link_select_t link_speed,

    output logic tmp_rxdv,
    output logic [7:0] tmp_rxd,
    output logic tmp_rxerr
);
// input DDR buffers =======================================================================
logic _rxdv, _rxerr;
logic [7:0] _rxd;

altddio_in #( /* RX enable and data capture */
  .intended_device_family("Cyclone V"),
  .invert_input_clocks("OFF"),
  .lpm_hint("UNUSED"),
  .lpm_type("altddio_in"),
  .power_up_high("OFF"),
  .width(5)
) rxio (
  .inclock(~eth_rxclk),
  .datain({eth_rxdv, eth_rxd}),
  .dataout_h({_rxerr, _rxd[7:4]}),
  .dataout_l({_rxdv, _rxd[3:0]}),
  .aclr(1'b0),
  .aset(1'b0),
  .inclocken(1'b1),
  .sclr(1'b0),
  .sset(1'b0)
);

assign tmp_rxdv = _rxdv;
assign tmp_rxd = _rxd;
assign tmp_rxerr = _rxerr;

// input synchronizer =======================================================================
logic rxdv_sync, rxerr_sync;
logic [7:0] rxd_sync;

vector_fifo_sync #(
  .pWIDTH(9)
) mii_sync_rx (
  .link_speed(link_speed),
  .clock_in(eth_rxclk),
  .ivalid(_rxdv),
  .ivector({_rxerr, _rxd}),
  .clock_out(clk),
  .ovalid(rxdv_sync),
  .ovector({rxerr_sync, rxd_sync})
);

// output DDR buffers =======================================================================
logic txen_d; /* Transmit enable signal */
logic [7:0] txd_d; // transmit data signal

assign eth_txclk = eth_txclk_phy; /* ToDo: Try to get rid of it */

wire txerr = txen_d ^ mii_tx.tx_error;

altddio_out #( // TX data generation
  .extend_oe_disable("OFF"),
  .intended_device_family("Cyclone V"),
  .invert_output("OFF"),
  .lpm_hint("UNUSED"),
  .lpm_type("altddio_out"),
  .oe_reg("UNREGISTERED"),
  .power_up_high("OFF"),
  .width(5)
) txio (
  .datain_h({txen_d, txd_d[3:0]}),
  .datain_l({txerr, txd_d[7:4]}),
  .outclock(eth_txck_in),
  .dataout({eth_txdv, eth_txd}),
  .aclr(1'b0),
  .aset(1'b0),
  .oe(1'b1),
  .oe_out(),
  .outclocken(1'b1),
  .sclr(1'b0),
  .sset(1'b0)
);
//==========================================================================================
logic [31:0] rx_crc, tx_crc;

function [31:0] crc_table;
input [3:0] addr;
  case (addr)
    0: crc_table = 32'h4DBDF21C;
    1: crc_table = 32'h500AE278;
    2: crc_table = 32'h76D3D2D4;
    3: crc_table = 32'h6B64C2B0;
    4: crc_table = 32'h3B61B38C;
    5: crc_table = 32'h26D6A3E8;
    6: crc_table = 32'h000F9344;
    7: crc_table = 32'h1DB88320;
    8: crc_table = 32'hA005713C;
    9: crc_table = 32'hBDB26158;
    10: crc_table = 32'h9B6B51F4;
    11: crc_table = 32'h86DC4190;
    12: crc_table = 32'hD6D930AC;
    13: crc_table = 32'hCB6E20C8;
    14: crc_table = 32'hEDB71064;
    default: crc_table = 32'hF0000000;
  endcase
endfunction

logic [31:0] rx_crc1, rx_crc2;
assign rx_crc1 = rx_crc[31:4] ^ crc_table(
  rx_crc[3:0] ^ rxd[3:0]
),
rx_crc2 = rx_crc1[31:4] ^ crc_table(
  rx_crc1[3:0] ^ rxd[7:4]
);

logic [31:0] tx_crc1, tx_crc2;
assign tx_crc1 = tx_crc[31:4] ^ crc_table(tx_crc[3:0] ^ mii_tx.data_tx[3:0]);
assign tx_crc2 = tx_crc1[31:4] ^ crc_table(tx_crc1[3:0] ^ mii_tx.data_tx[7:4]);

//==========================================================================================
logic [2 : 0] rx_pre_en;
logic valid_frame;
logic rxdv, rxdv_del;
logic [7 : 0] rxd;
logic rx_ff;
logic preamb_err_flg, min_frame_err_flg;
logic [3 : 0] min_length_cnt;
logic [7 : 0] link_cnt;
logic valid_rx_link;
logic str_100;

//assign rx_stat.line_err = (rx_stat.rx_fl & rxdv) | preamb_err_flg;

assign valid_rx = valid_rx_link && str_100;

always_ff @(posedge clk) begin : RX_MII_PROCESS
  if (~rst_n) begin
    rxdv <= 'd0;
    rxd <= 'd0;
    rxdv_del <= 'd0;
    rx_pre_en <= 'd0;
    rx_stat.rx_fl <= 'd0;
    rx_stat.crc_val <= 'd0;
    rx_stat.line_err = 'd0;
    valid_frame <= 'd0;
    preamb_err_flg <= 'd1;
    min_frame_err_flg <= 1'd1;
    min_length_cnt <= 'd0;
    valid_rx_link <= 'd0;
    data_rx <= 'd0;
    link_cnt <= 'd0;
    rx_ff <= 'd0;
    str_100 <= 'd0;
  end
  else begin
    rxdv_del <= rxdv;

    if (link_speed == LINK_1000) begin
      rxdv <= rxdv_sync;
      rxd <= rxd_sync;
      rx_ff <= 1'd1;
      str_100 <= 1'd1;
      link_cnt <= 'd0;
    end
    else begin
      rxdv <= rxdv_sync;
      str_100 <= rxdv & rx_ff;
      if (rxdv_sync)
        rxd <= {rxd_sync[7:4], rxd[7:4]};
      if (rxdv) begin
        if (link_speed == LINK_100)
          link_cnt <= 'd15;
        else
          link_cnt <= 'd150;
        rx_ff <= ~rx_ff;
      end
      else if (|link_cnt)
        link_cnt <= link_cnt - 1'd1;
      else
        rx_ff <= 'd0;
    end

    data_rx <= rxd;

    /* ABI: If we set valid_rx_link we must set rx_stat.rx_fl in the end. And vice versa! */
    if (rxdv & rx_ff) begin // data valid from mii
      rx_stat.rx_fl <= 'd0;
      rx_stat.crc_val <= 'd0;
      rx_stat.line_err = 'd0;
      valid_rx_link <= valid_frame;

      if (valid_frame) begin
        rx_crc <= rx_crc2;
        if (~&min_length_cnt)
          min_length_cnt <= min_length_cnt + 1'd1;
        else
          min_frame_err_flg <= 'd0;
      end
      else begin
        if (rxd == 8'h55)
          rx_pre_en <= rx_pre_en + 'd1;
        else
          rx_pre_en <= 'd0;

        if ((rx_pre_en == 3'd7) & (rxd == 8'hD5)) begin
          valid_frame <= 1'd1;
          rx_crc <= 'd0;
          preamb_err_flg <= 'd0;
          min_length_cnt <= 'd0;
        end
      end
    end
    else if (((link_speed == LINK_1000) && rxdv_del) || (link_speed != LINK_1000) && (link_cnt == 'd1)) begin
      rx_stat.rx_fl <= valid_rx_link;
      if (preamb_err_flg || min_frame_err_flg) begin
        rx_stat.crc_val <= 'd0;
        rx_stat.line_err = 1'd1;
      end
      else if (valid_rx_link) begin
        rx_stat.crc_val <= (rx_crc == 32'h2144DF1C);
        rx_stat.line_err = 'd0;
      end
      else begin
        rx_stat.crc_val <= 'd0;
        rx_stat.line_err = 1'd1;
      end

      valid_rx_link <= 'd0;
      valid_frame  <= 'd0;
      rx_pre_en <= 'd0;
      preamb_err_flg <= 'd1;
      min_length_cnt <= 'd0;
      min_frame_err_flg <= 1'd1;
    end
    else if (link_cnt == 'd0) begin
      rx_pre_en <= 'd0;
      rx_stat.rx_fl <= 'd0;
      rx_stat.crc_val <= 'd0;
      rx_stat.line_err = 'd0;
      valid_frame <= 'd0;
      preamb_err_flg <= 'd1;
      min_length_cnt <= 'd0;
      min_frame_err_flg <= 1'd1;
      valid_rx_link <= 'd0;
    end
  end
end
//==========================================================================================
logic [31:0] tx_pack_crc;
logic tx_crc_set;
logic [7:0] data_tx_del, data_tx_del_1G;
logic valid_tx_del, valid_tx_del_1G;
logic [2:0] tx_cnt;
logic tx_crc_en, tx_crc_en_1G;

delay_chain #( // forming preambule strobe
  .width(8 + 1),
  .depth(8)
) dc_tx (
  eth_txck_in,
  {mii_tx.valid_tx, mii_tx.data_tx},
  {valid_tx_del_1G, data_tx_del_1G}
);

delay_chain #(
  .depth(4)
) dc_tx_crc (
  eth_txck_in,
  valid_tx_del_1G,
  tx_crc_en_1G
);

assign valid_tx_del = valid_tx_del_1G;
assign data_tx_del = data_tx_del_1G;
assign tx_crc_en = tx_crc_en_1G;

function [7:0] byteselect(input [31:0] d, input [1:0] i); // byte select from the word
  case (i)
    2'd3: byteselect = d[31:24];
    2'd2: byteselect = d[23:16];
    2'd1: byteselect = d[15:8];
    default: byteselect = d[7:0];
  endcase
endfunction
wire [7:0] bs_res = byteselect(tx_pack_crc, tx_cnt[1:0]);

// 1Gbit/s, eth_txck_in = 125 MHz
// 100Mbit/s, eth_txck_in = 12.5 MHz
// 10Mbit/s, eth_txck_in = 1.25 MHz
always_ff @(posedge eth_txck_in) begin : TX_MII_PROCESS
  if (~rst_n) begin
    txd_d <= 'd0;
    txen_d <= 'd0;
  end
  else begin
    if (mii_tx.valid_tx) begin
      tx_crc <= tx_crc2;
      tx_crc_set <= 1'd1;
    end
    else begin
      tx_crc_set <= 1'd0;
      tx_crc <= 'd0;
      if (tx_crc_set)
        tx_pack_crc <= tx_crc;
    end

    txen_d <= mii_tx.valid_tx | tx_crc_en;

    if (~valid_tx_del & tx_crc_en) begin
      txd_d  <= bs_res;
      tx_cnt <= tx_cnt + 1'd1;
    end
    else if (valid_tx_del) begin
      txd_d <= data_tx_del;
      tx_cnt <= 'd0;
    end
    else if (mii_tx.valid_tx) begin
      tx_cnt <= tx_cnt - 1'd1;
      if (tx_cnt == 'd0)
        txd_d <= 8'hD5;
      else
        txd_d <= 8'h55;
    end
    else begin
      tx_cnt <= 3'd7;
      txd_d <= 'd0;
    end
  end
end

endmodule
